//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Departmen;t                                              --
//-------------------------------------------------------------------------


module boxhead( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK,     //SDRAM Clock
             //Audio
			 input	AUD_ADCDAT,
			 input AUD_DACLRCK,
			 input AUD_ADCLRCK,
			 input AUD_BCLK,
			 output logic AUD_DACDAT,
			 output logic AUD_XCK,
			 output logic I2C_SCLK,
			 output logic I2C_SDAT
                    );
    
    logic Reset_h, Clk;
    logic [7:0] keycode;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            .from_sw_reset(hpi_reset),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),
                            .OTG_RST_N(OTG_RST_N)
    );
     
     nios_system nios_system(
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
                             .otg_hpi_reset_export(hpi_reset)
    );
    
    // Audio Part
    // INIT: input logic for interface, generated by audio.
    // INIT_FINSH: Output logic for interface.
    // data_over: sample sync pulse
    logic INIT_FINISH, data_over, INIT;
    // Add is the pointer to the memory of target audio.
	logic [16:0] Add;
    // output audio signal, to the interface to play
	logic [16:0] music_content;
    logic[16:0] music_frequency;
    always_comb begin
		music_frequency = 16'd84;
	end
    audio audio1 (.*, .Reset(Reset_h));
	music music1 (.*);
    audio_interface music_int ( .LDATA(music_content), 
								.RDATA(music_content),
								.CLK(Clk),
								.Reset(Reset_h), 
								.INIT(INIT),
								.INIT_FINISH(INIT_FINISH),
								.adc_full(adc_full),
								.data_over(data_over),
								.AUD_MCLK(AUD_XCK),
								.AUD_BCLK(AUD_BCLK),     
								.AUD_ADCDAT(AUD_ADCDAT),
								.AUD_DACDAT(AUD_DACDAT),
								.AUD_DACLRCK(AUD_DACLRCK),
								.AUD_ADCLRCK(AUD_ADCLRCK),
								.I2C_SDAT(I2C_SDAT),
								.I2C_SCLK(I2C_SCLK),
								.ADCDATA(ADCDATA),
	);
    // VGA part
    logic [9:0] DrawX, DrawY;
    logic [8:0] PixelX, PixelY;

    logic [31:0] bkg_address;
    logic [15:0] player_address;
    logic [4:0] bkg_index;
    logic [4:0] player_index;
    logic [23:0] bkg_color;
    logic [23:0] player_color;

    logic is_player;

    assign PixelX = DrawX[9:1];
    assign PixelY = DrawY[9:1];

    assign bkg_address = PixelX + PixelY * 320;

    vga_controller vga_controller_inst(
        .*,
        .Reset(Reset_h),
        .hs(VGA_HS),
        .vs(VGA_VS),
        .pixel_clk(VGA_CLK),
        .blank(VGA_BLANK_N),
        .sync(VGA_SYNC_N)
    );

    backgroundRAM background_ram(
        .*,
        .data_In(),
        .write_address(),
        .read_address(bkg_address),
        .we(),
        .data_Out(bkg_index)
    );

    player player_inst(
        .*,
        .Reset(Reset_h),
        .frame_clk(VGA_VS),
        .keycode(keycode),
        .is_obj(is_player),
        .Obj_address(player_address)
    );

    playerROM playerROM_inst(
        .Clk(Clk),
        .read_address(player_address),
        .data_Out(player_index)
    );

    palette bkg_palette_inst(
        .*,
        .read_address(bkg_index),
        .data_Out(bkg_color)
    );

    palette player_palette_inst(
        .*,
        .read_address(player_index),
        .data_Out(player_color)
    );

    always_comb begin
        // If background is player and it's not red(sprite background color)
        if((is_player == 1'b1) && (player_index != 5'h0)) begin
            VGA_R = player_color[23:16];
            VGA_G = player_color[15:8];
            VGA_B = player_color[7:0];
        end
        else begin
            VGA_R = bkg_color[23:16];
            VGA_G = bkg_color[15:8];
            VGA_B = bkg_color[7:0];
        end

    end

    assign HEX0 = 7'hFF;
    assign HEX1 = 7'hFF; 

    // Display keycode on hex display
    // HexDriver hex_inst_0 (keycode[3:0], HEX0);
    // HexDriver hex_inst_1 (keycode[7:4], HEX1);

    
endmodule
